-- FC Package --

-- high-speed/low-power group
-- Fiore, Neri, Zheng
-- 
-- keyword in MAIUSCOLO (es: STD_LOGIC)
-- dati in minuscolo (es: data_in)
-- segnali di controllo in MAIUSCOLO (es: EN)
-- componenti instanziati con l'iniziale maiuscola (es: Shift_register_1)
-- i segnali attivi bassi con _n finale (es: RST_n)

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;


package FC_struct_pkg is

	CONSTANT INPUT_NEURONS_FC1   	: POSITIVE := 400;
	CONSTANT OUTPUT_NEURONS_FC1   : POSITIVE := 120;
	
	CONSTANT INPUT_NEURONS_FC2   	: POSITIVE := 120;
	CONSTANT OUTPUT_NEURONS_FC2   : POSITIVE := 84;
	
	CONSTANT INPUT_NEURONS_FC3   	: POSITIVE := 84;
	CONSTANT OUTPUT_NEURONS_FC3   : POSITIVE := 10;

	CONSTANT BIAS_SIZE      	: POSITIVE := 8;	
	CONSTANT WEIGHT_SIZE    	: POSITIVE := 8;
	CONSTANT OUTPUT_SIZE 		: POSITIVE := 8;
	CONSTANT INPUT_SIZE    		: POSITIVE := 8;
	
	CONSTANT N_MAC_FC1			: POSITIVE := 24;
	CONSTANT N_MAC_FC2			: POSITIVE := 21;
	CONSTANT N_MAC_FC3			: POSITIVE := 10;
	
	CONSTANT EXTRA_BIT			: NATURAL := 0;
	CONSTANT N_CYCLES_FC1		: POSITIVE :=5;
	CONSTANT N_CYCLES_FC2		: POSITIVE :=4;
	
	CONSTANT SEL_MUX_IN_SIZE_FC1   : POSITIVE := 9; -- Parallelism of selector ( ceil(log2(INPUT_NEURONS)) )
	CONSTANT SEL_MUX_IN_SIZE_FC2   : POSITIVE := 7; -- Parallelism of selector ( ceil(log2(INPUT_NEURONS)) )
	CONSTANT SEL_MUX_IN_SIZE_FC3   : POSITIVE := 7; -- Parallelism of selector ( ceil(log2(INPUT_NEURONS)) )
	
	TYPE weights_struct_FC1 IS ARRAY(N_MAC_FC1-1 DOWNTO 0) of STD_LOGIC_VECTOR(WEIGHT_SIZE-1 DOWNTO 0);
	TYPE weights_struct_FC2 IS ARRAY(N_MAC_FC2-1 DOWNTO 0) of STD_LOGIC_VECTOR(WEIGHT_SIZE-1 DOWNTO 0);
	TYPE weights_struct_FC3 IS ARRAY(N_MAC_FC3-1 DOWNTO 0) of STD_LOGIC_VECTOR(WEIGHT_SIZE-1 DOWNTO 0);
	
	TYPE bias_struct_FC1 IS ARRAY(N_MAC_FC1-1 DOWNTO 0) OF STD_LOGIC_VECTOR(BIAS_SIZE-1 DOWNTO 0);
	TYPE bias_struct_FC2 IS ARRAY(N_MAC_FC2-1 DOWNTO 0) OF STD_LOGIC_VECTOR(BIAS_SIZE-1 DOWNTO 0);
	TYPE bias_struct_FC3 IS ARRAY(N_MAC_FC3-1 DOWNTO 0) OF STD_LOGIC_VECTOR(BIAS_SIZE-1 DOWNTO 0);
	
	TYPE bias_mac_struct_FC1 IS ARRAY(N_MAC_FC1-1 DOWNTO 0) OF STD_LOGIC_VECTOR(2*BIAS_SIZE+EXTRA_BIT-2 DOWNTO 0);
	TYPE bias_mac_struct_FC2 IS ARRAY(N_MAC_FC2-1 DOWNTO 0) OF STD_LOGIC_VECTOR(2*BIAS_SIZE+EXTRA_BIT-2 DOWNTO 0);
	TYPE bias_mac_struct_FC3 IS ARRAY(N_MAC_FC3-1 DOWNTO 0) OF STD_LOGIC_VECTOR(2*BIAS_SIZE+EXTRA_BIT-2 DOWNTO 0);
	
	TYPE out_from_mac_FC1 IS ARRAY(N_MAC_FC1-1 DOWNTO 0) OF STD_LOGIC_VECTOR(OUTPUT_SIZE-1 DOWNTO 0);
	TYPE out_from_mac_FC2 IS ARRAY(N_MAC_FC2-1 DOWNTO 0) OF STD_LOGIC_VECTOR(OUTPUT_SIZE-1 DOWNTO 0);
	TYPE out_from_mac_FC3 IS ARRAY(N_MAC_FC3-1 DOWNTO 0) OF STD_LOGIC_VECTOR(OUTPUT_SIZE-1 DOWNTO 0);
	
end package;