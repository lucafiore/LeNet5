library verilog;
use verilog.vl_types.all;
entity seq_SDFFS_X2 is
    // This module cannot be connected to from
    // VHDL because it has unnamed ports.
end seq_SDFFS_X2;
